module AnalogToUInt (a, b);
  inout [0:0] a;
  output [0:0] b;
  assign b = a;
endmodule
